netcdf exampl2 {
dimensions:
	Time = UNLIMITED ; // (1 currently)
	DateStrLen = 19 ;
	west_east = 429 ;
	south_north = 468 ;
	num_press_levels_stag = 11 ;
variables:
	char Times(Time, DateStrLen) ;
	float XLAT(Time, south_north, west_east) ;
		XLAT:FieldType = 104 ;
		XLAT:MemoryOrder = "XY " ;
		XLAT:description = "LATITUDE, SOUTH IS NEGATIVE" ;
		XLAT:units = "degree_north" ;
		XLAT:stagger = "" ;
		XLAT:coordinates = "XLONG XLAT" ;
	float XLONG(Time, south_north, west_east) ;
		XLONG:FieldType = 104 ;
		XLONG:MemoryOrder = "XY " ;
		XLONG:description = "LONGITUDE, WEST IS NEGATIVE" ;
		XLONG:units = "degree_east" ;
		XLONG:stagger = "" ;
		XLONG:coordinates = "XLONG XLAT" ;
	float Q2(Time, south_north, west_east) ;
		Q2:FieldType = 104 ;
		Q2:MemoryOrder = "XY " ;
		Q2:description = "QV at 2 M" ;
		Q2:units = "kg kg-1" ;
		Q2:stagger = "" ;
		Q2:coordinates = "XLONG XLAT XTIME" ;
	float T2(Time, south_north, west_east) ;
		T2:FieldType = 104 ;
		T2:MemoryOrder = "XY " ;
		T2:description = "TEMP at 2 M" ;
		T2:units = "K" ;
		T2:stagger = "" ;
		T2:coordinates = "XLONG XLAT XTIME" ;
	float TH2(Time, south_north, west_east) ;
		TH2:FieldType = 104 ;
		TH2:MemoryOrder = "XY " ;
		TH2:description = "POT TEMP at 2 M" ;
		TH2:units = "K" ;
		TH2:stagger = "" ;
		TH2:coordinates = "XLONG XLAT XTIME" ;
	float PSFC(Time, south_north, west_east) ;
		PSFC:FieldType = 104 ;
		PSFC:MemoryOrder = "XY " ;
		PSFC:description = "SFC PRESSURE" ;
		PSFC:units = "Pa" ;
		PSFC:stagger = "" ;
		PSFC:coordinates = "XLONG XLAT XTIME" ;
	float U10(Time, south_north, west_east) ;
		U10:FieldType = 104 ;
		U10:MemoryOrder = "XY " ;
		U10:description = "U at 10 M" ;
		U10:units = "m s-1" ;
		U10:stagger = "" ;
		U10:coordinates = "XLONG XLAT XTIME" ;
	float V10(Time, south_north, west_east) ;
		V10:FieldType = 104 ;
		V10:MemoryOrder = "XY " ;
		V10:description = "V at 10 M" ;
		V10:units = "m s-1" ;
		V10:stagger = "" ;
		V10:coordinates = "XLONG XLAT XTIME" ;
	float LPI(Time, south_north, west_east) ;
		LPI:FieldType = 104 ;
		LPI:MemoryOrder = "XY " ;
		LPI:description = "Lightning Potential Index" ;
		LPI:units = "m^2 s-2" ;
		LPI:stagger = "" ;
		LPI:coordinates = "XLONG XLAT XTIME" ;
	float ACSNOW(Time, south_north, west_east) ;
		ACSNOW:FieldType = 104 ;
		ACSNOW:MemoryOrder = "XY " ;
		ACSNOW:description = "ACCUMULATED SNOW" ;
		ACSNOW:units = "kg m-2" ;
		ACSNOW:stagger = "" ;
		ACSNOW:coordinates = "XLONG XLAT XTIME" ;
	float RAINC(Time, south_north, west_east) ;
		RAINC:FieldType = 104 ;
		RAINC:MemoryOrder = "XY " ;
		RAINC:description = "ACCUMULATED TOTAL CUMULUS PRECIPITATION" ;
		RAINC:units = "mm" ;
		RAINC:stagger = "" ;
		RAINC:coordinates = "XLONG XLAT XTIME" ;
	float RAINNC(Time, south_north, west_east) ;
		RAINNC:FieldType = 104 ;
		RAINNC:MemoryOrder = "XY " ;
		RAINNC:description = "ACCUMULATED TOTAL GRID SCALE PRECIPITATION" ;
		RAINNC:units = "mm" ;
		RAINNC:stagger = "" ;
		RAINNC:coordinates = "XLONG XLAT XTIME" ;
	float SNOWNC(Time, south_north, west_east) ;
		SNOWNC:FieldType = 104 ;
		SNOWNC:MemoryOrder = "XY " ;
		SNOWNC:description = "ACCUMULATED TOTAL GRID SCALE SNOW AND ICE" ;
		SNOWNC:units = "mm" ;
		SNOWNC:stagger = "" ;
		SNOWNC:coordinates = "XLONG XLAT XTIME" ;
	float GRAUPELNC(Time, south_north, west_east) ;
		GRAUPELNC:FieldType = 104 ;
		GRAUPELNC:MemoryOrder = "XY " ;
		GRAUPELNC:description = "ACCUMULATED TOTAL GRID SCALE GRAUPEL" ;
		GRAUPELNC:units = "mm" ;
		GRAUPELNC:stagger = "" ;
		GRAUPELNC:coordinates = "XLONG XLAT XTIME" ;
	float HAILNC(Time, south_north, west_east) ;
		HAILNC:FieldType = 104 ;
		HAILNC:MemoryOrder = "XY " ;
		HAILNC:description = "ACCUMULATED TOTAL GRID SCALE HAIL" ;
		HAILNC:units = "mm" ;
		HAILNC:stagger = "" ;
		HAILNC:coordinates = "XLONG XLAT XTIME" ;
	float SWDOWN(Time, south_north, west_east) ;
		SWDOWN:FieldType = 104 ;
		SWDOWN:MemoryOrder = "XY " ;
		SWDOWN:description = "DOWNWARD SHORT WAVE FLUX AT GROUND SURFACE" ;
		SWDOWN:units = "W m-2" ;
		SWDOWN:stagger = "" ;
		SWDOWN:coordinates = "XLONG XLAT XTIME" ;
	float SWDOWNC(Time, south_north, west_east) ;
		SWDOWNC:FieldType = 104 ;
		SWDOWNC:MemoryOrder = "XY " ;
		SWDOWNC:description = "DOWNWARD CLEAR-SKY SHORT WAVE FLUX AT GROUND SURFACE" ;
		SWDOWNC:units = "W m-2" ;
		SWDOWNC:stagger = "" ;
		SWDOWNC:coordinates = "XLONG XLAT XTIME" ;
	float PBLH(Time, south_north, west_east) ;
		PBLH:FieldType = 104 ;
		PBLH:MemoryOrder = "XY " ;
		PBLH:description = "PBL HEIGHT" ;
		PBLH:units = "m" ;
		PBLH:stagger = "" ;
		PBLH:coordinates = "XLONG XLAT XTIME" ;
	float HFX(Time, south_north, west_east) ;
		HFX:FieldType = 104 ;
		HFX:MemoryOrder = "XY " ;
		HFX:description = "UPWARD HEAT FLUX AT THE SURFACE" ;
		HFX:units = "W m-2" ;
		HFX:stagger = "" ;
		HFX:coordinates = "XLONG XLAT XTIME" ;
	float QFX(Time, south_north, west_east) ;
		QFX:FieldType = 104 ;
		QFX:MemoryOrder = "XY " ;
		QFX:description = "UPWARD MOISTURE FLUX AT THE SURFACE" ;
		QFX:units = "kg m-2 s-1" ;
		QFX:stagger = "" ;
		QFX:coordinates = "XLONG XLAT XTIME" ;
	float LH(Time, south_north, west_east) ;
		LH:FieldType = 104 ;
		LH:MemoryOrder = "XY " ;
		LH:description = "LATENT HEAT FLUX AT THE SURFACE" ;
		LH:units = "W m-2" ;
		LH:stagger = "" ;
		LH:coordinates = "XLONG XLAT XTIME" ;
	float WSPD10MAX(Time, south_north, west_east) ;
		WSPD10MAX:FieldType = 104 ;
		WSPD10MAX:MemoryOrder = "XY " ;
		WSPD10MAX:description = "WIND SPD MAX 10 M" ;
		WSPD10MAX:units = "m s-1" ;
		WSPD10MAX:stagger = "" ;
		WSPD10MAX:coordinates = "XLONG XLAT XTIME" ;
	float W_UP_MAX(Time, south_north, west_east) ;
		W_UP_MAX:FieldType = 104 ;
		W_UP_MAX:MemoryOrder = "XY " ;
		W_UP_MAX:description = "MAX Z-WIND UPDRAFT" ;
		W_UP_MAX:units = "m s-1" ;
		W_UP_MAX:stagger = "" ;
		W_UP_MAX:coordinates = "XLONG XLAT XTIME" ;
	float W_DN_MAX(Time, south_north, west_east) ;
		W_DN_MAX:FieldType = 104 ;
		W_DN_MAX:MemoryOrder = "XY " ;
		W_DN_MAX:description = "MAX Z-WIND DOWNDRAFT" ;
		W_DN_MAX:units = "m s-1" ;
		W_DN_MAX:stagger = "" ;
		W_DN_MAX:coordinates = "XLONG XLAT XTIME" ;
	float REFD_MAX(Time, south_north, west_east) ;
		REFD_MAX:FieldType = 104 ;
		REFD_MAX:MemoryOrder = "XY " ;
		REFD_MAX:description = "MAX DERIVED RADAR REFL" ;
		REFD_MAX:units = "dbZ" ;
		REFD_MAX:stagger = "" ;
		REFD_MAX:coordinates = "XLONG XLAT XTIME" ;
	float UP_HELI_MAX(Time, south_north, west_east) ;
		UP_HELI_MAX:FieldType = 104 ;
		UP_HELI_MAX:MemoryOrder = "XY " ;
		UP_HELI_MAX:description = "MAX UPDRAFT HELICITY" ;
		UP_HELI_MAX:units = "m2 s-2" ;
		UP_HELI_MAX:stagger = "" ;
		UP_HELI_MAX:coordinates = "XLONG XLAT XTIME" ;
	float W_MEAN(Time, south_north, west_east) ;
		W_MEAN:FieldType = 104 ;
		W_MEAN:MemoryOrder = "XY " ;
		W_MEAN:description = "HOURLY MEAN Z-WIND" ;
		W_MEAN:units = "m s-1" ;
		W_MEAN:stagger = "" ;
		W_MEAN:coordinates = "XLONG XLAT XTIME" ;
	float GRPL_MAX(Time, south_north, west_east) ;
		GRPL_MAX:FieldType = 104 ;
		GRPL_MAX:MemoryOrder = "XY " ;
		GRPL_MAX:description = "MAX COL INT GRAUPEL" ;
		GRPL_MAX:units = "kg m-2" ;
		GRPL_MAX:stagger = "" ;
		GRPL_MAX:coordinates = "XLONG XLAT XTIME" ;
	float UH(Time, south_north, west_east) ;
		UH:FieldType = 104 ;
		UH:MemoryOrder = "XY " ;
		UH:description = "UPDRAFT HELICITY" ;
		UH:units = "m2 s-2" ;
		UH:stagger = "" ;
		UH:coordinates = "XLONG XLAT XTIME" ;
	float HAIL_MAX2D(Time, south_north, west_east) ;
		HAIL_MAX2D:FieldType = 104 ;
		HAIL_MAX2D:MemoryOrder = "XY " ;
		HAIL_MAX2D:description = "MAX HAIL DIAMETER ENTIRE COLUMN" ;
		HAIL_MAX2D:units = "m" ;
		HAIL_MAX2D:stagger = "" ;
		HAIL_MAX2D:coordinates = "XLONG XLAT XTIME" ;
	float P_PL(Time, num_press_levels_stag) ;
		P_PL:FieldType = 104 ;
		P_PL:MemoryOrder = "Z  " ;
		P_PL:description = "Pressure level data, Pressure" ;
		P_PL:units = "Pa" ;
		P_PL:stagger = "Z" ;
	float U_PL(Time, num_press_levels_stag, south_north, west_east) ;
		U_PL:FieldType = 104 ;
		U_PL:MemoryOrder = "XYZ" ;
		U_PL:description = "Pressure level data, U wind" ;
		U_PL:units = "m s-1" ;
		U_PL:stagger = "Z" ;
		U_PL:coordinates = "XLONG XLAT XTIME" ;
	float V_PL(Time, num_press_levels_stag, south_north, west_east) ;
		V_PL:FieldType = 104 ;
		V_PL:MemoryOrder = "XYZ" ;
		V_PL:description = "Pressure level data, V wind" ;
		V_PL:units = "m s-1" ;
		V_PL:stagger = "Z" ;
		V_PL:coordinates = "XLONG XLAT XTIME" ;
	float T_PL(Time, num_press_levels_stag, south_north, west_east) ;
		T_PL:FieldType = 104 ;
		T_PL:MemoryOrder = "XYZ" ;
		T_PL:description = "Pressure level data, Temperature" ;
		T_PL:units = "K" ;
		T_PL:stagger = "Z" ;
		T_PL:coordinates = "XLONG XLAT XTIME" ;
	float RH_PL(Time, num_press_levels_stag, south_north, west_east) ;
		RH_PL:FieldType = 104 ;
		RH_PL:MemoryOrder = "XYZ" ;
		RH_PL:description = "Pressure level data, Relative humidity" ;
		RH_PL:units = "%" ;
		RH_PL:stagger = "Z" ;
		RH_PL:coordinates = "XLONG XLAT XTIME" ;
	float GHT_PL(Time, num_press_levels_stag, south_north, west_east) ;
		GHT_PL:FieldType = 104 ;
		GHT_PL:MemoryOrder = "XYZ" ;
		GHT_PL:description = "Pressure level data, Geopotential Height" ;
		GHT_PL:units = "m" ;
		GHT_PL:stagger = "Z" ;
		GHT_PL:coordinates = "XLONG XLAT XTIME" ;
	float S_PL(Time, num_press_levels_stag, south_north, west_east) ;
		S_PL:FieldType = 104 ;
		S_PL:MemoryOrder = "XYZ" ;
		S_PL:description = "Pressure level data, Speed" ;
		S_PL:units = "m s-1" ;
		S_PL:stagger = "Z" ;
		S_PL:coordinates = "XLONG XLAT XTIME" ;
	float TD_PL(Time, num_press_levels_stag, south_north, west_east) ;
		TD_PL:FieldType = 104 ;
		TD_PL:MemoryOrder = "XYZ" ;
		TD_PL:description = "Pressure level data, Dew point temperature" ;
		TD_PL:units = "K" ;
		TD_PL:stagger = "Z" ;
		TD_PL:coordinates = "XLONG XLAT XTIME" ;
	float Q_PL(Time, num_press_levels_stag, south_north, west_east) ;
		Q_PL:FieldType = 104 ;
		Q_PL:MemoryOrder = "XYZ" ;
		Q_PL:description = "Pressure level data, Mixing ratio" ;
		Q_PL:units = "kg/kg" ;
		Q_PL:stagger = "Z" ;
		Q_PL:coordinates = "XLONG XLAT XTIME" ;

// global attributes:
		:TITLE = " OUTPUT FROM WRF V3.8.1 MODEL" ;
		:START_DATE = "2021-12-13_00:00:00" ;
		:WEST-EAST_GRID_DIMENSION = 430 ;
		:SOUTH-NORTH_GRID_DIMENSION = 469 ;
		:BOTTOM-TOP_GRID_DIMENSION = 50 ;
		:DX = 2500.f ;
		:DY = 2500.f ;
		:P_LEV_MISSING = -999.f ;
		:GRIDTYPE = "C" ;
		:DIFF_OPT = 2 ;
		:KM_OPT = 2 ;
		:DAMP_OPT = 0 ;
		:DAMPCOEF = 0.2f ;
		:KHDIF = 0.f ;
		:KVDIF = 0.f ;
		:MP_PHYSICS = 6 ;
		:RA_LW_PHYSICS = 4 ;
		:RA_SW_PHYSICS = 4 ;
		:SF_SFCLAY_PHYSICS = 1 ;
		:SF_SURFACE_PHYSICS = 3 ;
		:BL_PBL_PHYSICS = 1 ;
		:CU_PHYSICS = 0 ;
		:SF_LAKE_PHYSICS = 0 ;
		:SURFACE_INPUT_SOURCE = 1 ;
		:SST_UPDATE = 0 ;
		:GRID_FDDA = 0 ;
		:GFDDA_INTERVAL_M = 0 ;
		:GFDDA_END_H = 0 ;
		:GRID_SFDDA = 0 ;
		:SGFDDA_INTERVAL_M = 0 ;
		:SGFDDA_END_H = 0 ;
		:HYPSOMETRIC_OPT = 2 ;
		:USE_THETA_M = 0 ;
		:WEST-EAST_PATCH_START_UNSTAG = 1 ;
		:WEST-EAST_PATCH_END_UNSTAG = 429 ;
		:WEST-EAST_PATCH_START_STAG = 1 ;
		:WEST-EAST_PATCH_END_STAG = 430 ;
		:SOUTH-NORTH_PATCH_START_UNSTAG = 1 ;
		:SOUTH-NORTH_PATCH_END_UNSTAG = 468 ;
		:SOUTH-NORTH_PATCH_START_STAG = 1 ;
		:SOUTH-NORTH_PATCH_END_STAG = 469 ;
		:BOTTOM-TOP_PATCH_START_UNSTAG = 1 ;
		:BOTTOM-TOP_PATCH_END_UNSTAG = 49 ;
		:BOTTOM-TOP_PATCH_START_STAG = 1 ;
		:BOTTOM-TOP_PATCH_END_STAG = 50 ;
		:GRID_ID = 3 ;
		:PARENT_ID = 2 ;
		:I_PARENT_START = 162 ;
		:J_PARENT_START = 79 ;
		:PARENT_GRID_RATIO = 3 ;
		:DT = 14.f ;
		:CEN_LAT = 42.14218f ;
		:CEN_LON = 12.03256f ;
		:TRUELAT1 = 47.f ;
		:TRUELAT2 = 0.f ;
		:MOAD_CEN_LAT = 47.f ;
		:STAND_LON = 15.f ;
		:POLE_LAT = 90.f ;
		:POLE_LON = 0.f ;
		:GMT = 0.f ;
		:JULYR = 2021 ;
		:JULDAY = 347 ;
		:MAP_PROJ = 3 ;
		:MAP_PROJ_CHAR = "Mercator" ;
		:MMINLU = "MODIFIED_IGBP_MODIS_NOAH" ;
		:NUM_LAND_CAT = 21 ;
		:ISWATER = 17 ;
		:ISLAKE = 21 ;
		:ISICE = 15 ;
		:ISURBAN = 13 ;
		:ISOILWATER = 14 ;
}
